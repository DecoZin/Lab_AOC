library ieee;
use ieee.std_logic_1164.all;

entity mux31 is
    generic (
        largura_dado : natural := 32
    );
    port (
        dado_ent_0, dado_ent_1, dado_ent_2 : in std_logic_vector((largura_dado - 1) downto 0);
        sele_ent                           : in std_logic_vector(1 downto 0);
        dado_sai                           : out std_logic_vector((largura_dado - 1) downto 0)
    );
end mux31;

architecture dataflow of mux31 is
begin
    with sele_ent select
        dado_sai <= dado_ent_0 when "00",
                    dado_ent_1 when "01",
                    dado_ent_2 when "10",
                    (others => '0') when others; 
end dataflow;
